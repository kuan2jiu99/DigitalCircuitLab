// Hexadecimal numbers
`define HEX_0 4'h0
`define HEX_1 4'h1
`define HEX_2 4'h2
`define HEX_3 4'h3
`define HEX_4 4'h4
`define HEX_5 4'h5
`define HEX_6 4'h6
`define HEX_7 4'h7
`define HEX_8 4'h8
`define HEX_9 4'h9
`define HEX_A 4'hA
`define HEX_B 4'hB
`define HEX_C 4'hC
`define HEX_D 4'hD
`define HEX_E 4'hE
`define HEX_F 4'hF

// Extend keys
`define EX 1'b1
`define NOT_EX 1'b0

module output_control (
last_change,  // last_change from KeyboardDecoder.v
key_num  // encoded keyboard number
    );
    
input [8:0] last_change;
output reg [3:0] key_num; // W: UP(0), S: DOWN(1), A: LEFT(2), D:RIGHT(3)

// Combinational Logic : Encoder
always @*
    case (last_change)
        {`NOT_EX, `HEX_1, `HEX_D} : key_num = 4'd0; // W: UP
        {`NOT_EX, `HEX_1, `HEX_B} : key_num = 4'd1; // S: DOWN
        {`NOT_EX, `HEX_1, `HEX_C} : key_num = 4'd2; // A: LEFT
        {`NOT_EX, `HEX_2, `HEX_3} : key_num = 4'd3; // D: RIGHT
        default : key_num = 4'd0;
        endcase
        
endmodule